module tpumac_tb();


    logic clk; 
    logic rst_n;
    logic WrEn;
    logic en;

    logic signed [BITS_AB-1:0] Ain,
    logic signed [BITS_AB-1:0] Bin,
    logic signed [BITS_C-1:0] Cin,

    logic reg signed [BITS_AB-1:0] Aout,   
    logic reg signed [BITS_AB-1:0] Bout,
    logic reg signed [BITS_C-1:0] Cout


endmodule 